
`define HWC_ROM1_OFF
`define HWC_RAMCART128
`define HWC_BRAM_8B
`define MUTE_VOL -8192