
`include "../hwc.sv"


`define USE_MDP
`define USE_MCD


//`define MCD_MUTE
//`define MCD_DSP_OFF

