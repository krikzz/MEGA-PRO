
`define HWC_ROM1_ON
`define HWC_RAMCART128
`define HWC_BRAM_16B
`define MUTE_VOL 0