

`define HWC_ROM1_ON
`define MUTE_VOL 0
