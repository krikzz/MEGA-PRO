
`include "../hwc.sv"


`define USE_MDP
//`define USE_MCD
//`define DSP_OFF
