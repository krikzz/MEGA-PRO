
`include "../hwc.sv"
