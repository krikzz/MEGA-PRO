
`include "../hwc.sv"

