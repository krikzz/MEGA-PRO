
`include "../hwc.sv"


`define USE_MCD
`define MCD_MASTER


//`define MCD_MUTE
//`define MCD_DSP_OFF
