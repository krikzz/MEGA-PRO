

`define HWC_ROM1_OFF
`define MUTE_VOL -8192

