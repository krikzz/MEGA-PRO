
`include "../hwc.sv"


//`define USE_SST_SMD
//`define USE_CHEATS
